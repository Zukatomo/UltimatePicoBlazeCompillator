library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
library unisim;
use unisim.vcomponents.all;
entity lcd_prg is
    Port (      addressA : in std_logic_vector(9 downto 0);
 addressB : in std_logic_vector(9 downto 0);
                instructionA : out std_logic_vector(17 downto 0);
  instructionB : out std_logic_vector(17 downto 0);
               clk : in std_logic);
    end lcd_prg;
architecture low_level_definition of lcd_prg is
attribute INIT_00 : string;
attribute INIT_01 : string;
attribute INIT_02 : string;
attribute INIT_03 : string;
attribute INIT_04 : string;
attribute INIT_05 : string;
attribute INIT_06 : string;
attribute INIT_07 : string;
attribute INIT_08 : string;
attribute INIT_09 : string;
attribute INIT_0A : string;
attribute INIT_0B : string;
attribute INIT_0C : string;
attribute INIT_0D : string;
attribute INIT_0E : string;
attribute INIT_0F : string;
attribute INIT_10 : string;
attribute INIT_11 : string;
attribute INIT_12 : string;
attribute INIT_13 : string;
attribute INIT_14 : string;
attribute INIT_15 : string;
attribute INIT_16 : string;
attribute INIT_17 : string;
attribute INIT_18 : string;
attribute INIT_19 : string;
attribute INIT_1A : string;
attribute INIT_1B : string;
attribute INIT_1C : string;
attribute INIT_1D : string;
attribute INIT_1E : string;
attribute INIT_1F : string;
attribute INIT_20 : string;
attribute INIT_21 : string;
attribute INIT_22 : string;
attribute INIT_23 : string;
attribute INIT_24 : string;
attribute INIT_25 : string;
attribute INIT_26 : string;
attribute INIT_27 : string;
attribute INIT_28 : string;
attribute INIT_29 : string;
attribute INIT_2A : string;
attribute INIT_2B : string;
attribute INIT_2C : string;
attribute INIT_2D : string;
attribute INIT_2E : string;
attribute INIT_2F : string;
attribute INIT_30 : string;
attribute INIT_31 : string;
attribute INIT_32 : string;
attribute INIT_33 : string;
attribute INIT_34 : string;
attribute INIT_35 : string;
attribute INIT_36 : string;
attribute INIT_37 : string;
attribute INIT_38 : string;
attribute INIT_39 : string;
attribute INIT_3A : string;
attribute INIT_3B : string;
attribute INIT_3C : string;
attribute INIT_3D : string;
attribute INIT_3E : string;
attribute INIT_3F : string;
attribute INITP_00 : string;
attribute INITP_01 : string;
attribute INITP_02 : string;
attribute INITP_03 : string;
attribute INITP_04 : string;
attribute INITP_05 : string;
attribute INITP_06 : string;
attribute INITP_07 : string;
attribute INIT_00 of ram_1024_x_18  : label is "CCFF0B0006000C00EF000F010A0F1180107009CC08010798050604C6CE800E00";
attribute INIT_01 of ram_1024_x_18  : label is "90F05FB00F070F00CE800E00503A4DFF500C4C118C01CFFE0F000044C171C070";
attribute INIT_02 of ram_1024_x_18  : label is "400ED6C0060F0DFFCE800E01010010905C30551013101200581C4B208B01A100";
attribute INIT_03 of ram_1024_x_18  : label is "400EA1008005C60150404600400ECFFE0F0110705837570054374100E100D0A0";
attribute INIT_04 of ram_1024_x_18  : label is "CC0100520C32A0005449C001004DA0005C442F014FFD0F07400ECFFE0F010D00";
attribute INIT_05 of ram_1024_x_18  : label is "A000CC01CC01CC010C03A0005458CC010C0BA0005453CC0100570CC8A000544E";
attribute INIT_06 of ram_1024_x_18  : label is "0C0EA0008C07B8004C3A8C300C0E0C0E0C0E0C0EA0008C07B8004C3A8C30AC0F";
attribute INIT_07 of ram_1024_x_18  : label is "8C07B8004C3A8C300C0E0C0E0C0E0C0EA0008C07B8004C3A8C300C0E0C0E0C0E";
attribute INIT_08 of ram_1024_x_18  : label is "4600400EA1008005C60150404600A000544ECC010052A000544ECC010052A000";
attribute INIT_09 of ram_1024_x_18  : label is "09CC08010798050604C6400EA1008005C60150404600400EA1008005C6015040";
attribute INIT_0A of ram_1024_x_18  : label is "0506EF000F010A0F1180107009CC08010798050604C6EF000F010A0F11801070";
attribute INIT_0B of ram_1024_x_18  : label is "050600AF0A0F1180107009CC08010798050600BF0A0F1180107009CC08010798";
attribute INIT_0C of ram_1024_x_18  : label is "A0008C07B8004C3A8C300C0E0C0E0C0E0C0E00B70A0F1180107009CC08010798";
attribute INIT_0D of ram_1024_x_18  : label is "B8004C3A8C300C0E0C0E0C0E0C0EA0008C07B8004C3A8C300C0E0C0E0C0E0C0E";
attribute INIT_0E of ram_1024_x_18  : label is "400EA1008005C60150404600A000544ECC010052A000544ECC010052A0008C07";
attribute INIT_0F of ram_1024_x_18  : label is "90F05FB00F070F00400EA1008005C60150404600400EA1008005C60150404600";
attribute INIT_10 of ram_1024_x_18  : label is "8C300C0E0C0E0C0E0C0E00B70A0F1180107009CC08010798581C4B208B01A100";
attribute INIT_11 of ram_1024_x_18  : label is "0C0E0C0E0C0EA0008C07B8004C3A8C300C0E0C0E0C0E0C0EA0008C07B8004C3A";
attribute INIT_12 of ram_1024_x_18  : label is "50404600A000544ECC010052A000544ECC010052A0008C07B8004C3A8C300C0E";
attribute INIT_13 of ram_1024_x_18  : label is "400EA1008005C60150404600400EA1008005C60150404600400EA1008005C601";
attribute INIT_14 of ram_1024_x_18  : label is "0C0E00B70A0F1180107009CC08010798581C4B208B01A10090F05FB00F070F00";
attribute INIT_15 of ram_1024_x_18  : label is "8C07B8004C3A8C300C0E0C0E0C0E0C0EA0008C07B8004C3A8C300C0E0C0E0C0E";
attribute INIT_16 of ram_1024_x_18  : label is "CC010052A000544ECC010052A0008C07B8004C3A8C300C0E0C0E0C0E0C0EA000";
attribute INIT_17 of ram_1024_x_18  : label is "50404600400EA1008005C60150404600400EA1008005C60150404600A000544E";
attribute INIT_18 of ram_1024_x_18  : label is "107009CC08010798581C4B208B01A10090F05FB00F070F00400EA1008005C601";
attribute INIT_19 of ram_1024_x_18  : label is "0C0E0C0E0C0E0C0EA0008C07B8004C3A8C300C0E0C0E0C0E0C0E00B70A0F1180";
attribute INIT_1A of ram_1024_x_18  : label is "CC010052A0008C07B8004C3A8C300C0E0C0E0C0E0C0EA0008C07B8004C3A8C30";
attribute INIT_1B of ram_1024_x_18  : label is "8005C60150404600400EA1008005C60150404600A000544ECC010052A000544E";
attribute INIT_1C of ram_1024_x_18  : label is "581C4B208B01A10090F05FB00F070F00400EA1008005C60150404600400EA100";
attribute INIT_1D of ram_1024_x_18  : label is "0C0EA0005449C001A0005449C001A0005449C001A0005449C001A0005449C001";
attribute INIT_1E of ram_1024_x_18  : label is "0C0EA0008C07B8004C3A8C300C0E0C0E0C0E0C0EA0008C07B8004C3A8C300C0E";
attribute INIT_1F of ram_1024_x_18  : label is "A000544ECC010052A000544ECC010052A0008C07B8004C3A8C300C0E0C0E0C0E";
attribute INIT_20 of ram_1024_x_18  : label is "8005C60150404600400EA1008005C60150404600400EA1008005C60150404600";
attribute INIT_21 of ram_1024_x_18  : label is "8C07B8004C3A8C300C0E0C0E581C4B208B01A10090F05FB00F070F00400EA100";
attribute INIT_22 of ram_1024_x_18  : label is "4C3A8C300C0E0C0E0C0E0C0EA0008C07B8004C3A8C300C0E0C0E0C0E0C0EA000";
attribute INIT_23 of ram_1024_x_18  : label is "A1008005C60150404600A000544ECC010052A000544ECC010052A0008C07B800";
attribute INIT_24 of ram_1024_x_18  : label is "5FB00F070F00400EA1008005C60150404600400EA1008005C60150404600400E";
attribute INIT_25 of ram_1024_x_18  : label is "0C0E0C0E0C0E0C0EA0008C07B8004C3A8C300C0E0C0E581C4B208B01A10090F0";
attribute INIT_26 of ram_1024_x_18  : label is "CC010052A0008C07B8004C3A8C300C0E0C0E0C0E0C0EA0008C07B8004C3A8C30";
attribute INIT_27 of ram_1024_x_18  : label is "8005C60150404600400EA1008005C60150404600A000544ECC010052A000544E";
attribute INIT_28 of ram_1024_x_18  : label is "581C4B208B01A10090F05FB00F070F00400EA1008005C60150404600400EA100";
attribute INIT_29 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_2A of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_2B of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_2C of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_2D of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_2E of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_2F of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_30 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_31 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_32 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_33 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_34 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_35 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_36 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_37 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_38 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_39 of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_3A of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_3B of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_3C of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_3D of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_3E of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INIT_3F of ram_1024_x_18  : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INITP_00 of ram_1024_x_18 : label is "65AA996AA65AA994952D2DCB72DED2E0D5DE0DD5D080D0D5488DD63A80800008";
attribute INITP_01 of ram_1024_x_18 : label is "48D5DD5DD5DB7B7996AA65AA996AB0003000300020000200003577577576DEDE";
attribute INITP_02 of ram_1024_x_18 : label is "DD5DD5DB7B7996AA65AA996AB000D548D5DD5DD5DB7B7996AA65AA996AB000D5";
attribute INITP_03 of ram_1024_x_18 : label is "B7B7996AA65AA996ADB6DB6DD548D5DD5DD5DB7B7996AA65AA996AB000D548D5";
attribute INITP_04 of ram_1024_x_18 : label is "5DD5DB7B7996AA65AA996B5523577577576DEDE65AA996AA65AD548D5DD5DD5D";
attribute INITP_05 of ram_1024_x_18 : label is "00000000000000000000000000000000000000000000000000000000D548D5DD";
attribute INITP_06 of ram_1024_x_18 : label is "0000000000000000000000000000000000000000000000000000000000000000";
attribute INITP_07 of ram_1024_x_18 : label is "0000000000000000000000000000000000000000000000000000000000000000";
begin
--
  --Instantiate the Xilinx primitive for a block RAM
  ram_1024_x_18: RAMB16_S18
  --synthesis translate_off
  --INIT values repeated to define contents for functional simulation
generic map ( INIT_00 => X"CCFF0B0006000C00EF000F010A0F1180107009CC08010798050604C6CE800E00",
			  INIT_01 => X"90F05FB00F070F00CE800E00503A4DFF500C4C118C01CFFE0F000044C171C070",
			  INIT_02 => X"400ED6C0060F0DFFCE800E01010010905C30551013101200581C4B208B01A100",
			  INIT_03 => X"400EA1008005C60150404600400ECFFE0F0110705837570054374100E100D0A0",
			  INIT_04 => X"CC0100520C32A0005449C001004DA0005C442F014FFD0F07400ECFFE0F010D00",
			  INIT_05 => X"A000CC01CC01CC010C03A0005458CC010C0BA0005453CC0100570CC8A000544E",
			  INIT_06 => X"0C0EA0008C07B8004C3A8C300C0E0C0E0C0E0C0EA0008C07B8004C3A8C30AC0F",
			  INIT_07 => X"8C07B8004C3A8C300C0E0C0E0C0E0C0EA0008C07B8004C3A8C300C0E0C0E0C0E",
			  INIT_08 => X"4600400EA1008005C60150404600A000544ECC010052A000544ECC010052A000",
			  INIT_09 => X"09CC08010798050604C6400EA1008005C60150404600400EA1008005C6015040",
			  INIT_0A => X"0506EF000F010A0F1180107009CC08010798050604C6EF000F010A0F11801070",
			  INIT_0B => X"050600AF0A0F1180107009CC08010798050600BF0A0F1180107009CC08010798",
			  INIT_0C => X"A0008C07B8004C3A8C300C0E0C0E0C0E0C0E00B70A0F1180107009CC08010798",
			  INIT_0D => X"B8004C3A8C300C0E0C0E0C0E0C0EA0008C07B8004C3A8C300C0E0C0E0C0E0C0E",
			  INIT_0E => X"400EA1008005C60150404600A000544ECC010052A000544ECC010052A0008C07",
			  INIT_0F => X"90F05FB00F070F00400EA1008005C60150404600400EA1008005C60150404600",
			  INIT_10 => X"8C300C0E0C0E0C0E0C0E00B70A0F1180107009CC08010798581C4B208B01A100",
			  INIT_11 => X"0C0E0C0E0C0EA0008C07B8004C3A8C300C0E0C0E0C0E0C0EA0008C07B8004C3A",
			  INIT_12 => X"50404600A000544ECC010052A000544ECC010052A0008C07B8004C3A8C300C0E",
			  INIT_13 => X"400EA1008005C60150404600400EA1008005C60150404600400EA1008005C601",
			  INIT_14 => X"0C0E00B70A0F1180107009CC08010798581C4B208B01A10090F05FB00F070F00",
			  INIT_15 => X"8C07B8004C3A8C300C0E0C0E0C0E0C0EA0008C07B8004C3A8C300C0E0C0E0C0E",
			  INIT_16 => X"CC010052A000544ECC010052A0008C07B8004C3A8C300C0E0C0E0C0E0C0EA000",
			  INIT_17 => X"50404600400EA1008005C60150404600400EA1008005C60150404600A000544E",
			  INIT_18 => X"107009CC08010798581C4B208B01A10090F05FB00F070F00400EA1008005C601",
			  INIT_19 => X"0C0E0C0E0C0E0C0EA0008C07B8004C3A8C300C0E0C0E0C0E0C0E00B70A0F1180",
			  INIT_1A => X"CC010052A0008C07B8004C3A8C300C0E0C0E0C0E0C0EA0008C07B8004C3A8C30",
			  INIT_1B => X"8005C60150404600400EA1008005C60150404600A000544ECC010052A000544E",
			  INIT_1C => X"581C4B208B01A10090F05FB00F070F00400EA1008005C60150404600400EA100",
			  INIT_1D => X"0C0EA0005449C001A0005449C001A0005449C001A0005449C001A0005449C001",
			  INIT_1E => X"0C0EA0008C07B8004C3A8C300C0E0C0E0C0E0C0EA0008C07B8004C3A8C300C0E",
			  INIT_1F => X"A000544ECC010052A000544ECC010052A0008C07B8004C3A8C300C0E0C0E0C0E",
			  INIT_20 => X"8005C60150404600400EA1008005C60150404600400EA1008005C60150404600",
			  INIT_21 => X"8C07B8004C3A8C300C0E0C0E581C4B208B01A10090F05FB00F070F00400EA100",
			  INIT_22 => X"4C3A8C300C0E0C0E0C0E0C0EA0008C07B8004C3A8C300C0E0C0E0C0E0C0EA000",
			  INIT_23 => X"A1008005C60150404600A000544ECC010052A000544ECC010052A0008C07B800",
			  INIT_24 => X"5FB00F070F00400EA1008005C60150404600400EA1008005C60150404600400E",
			  INIT_25 => X"0C0E0C0E0C0E0C0EA0008C07B8004C3A8C300C0E0C0E581C4B208B01A10090F0",
			  INIT_26 => X"CC010052A0008C07B8004C3A8C300C0E0C0E0C0E0C0EA0008C07B8004C3A8C30",
			  INIT_27 => X"8005C60150404600400EA1008005C60150404600A000544ECC010052A000544E",
			  INIT_28 => X"581C4B208B01A10090F05FB00F070F00400EA1008005C60150404600400EA100",
			  INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
			  INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
			  INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
			  INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
			  INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
			  INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
			  INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
			  INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
			  INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
			  INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
			  INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
			  INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
			  INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
			  INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
			  INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
			  INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
			  INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
			  INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
			  INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
			  INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
			  INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
			  INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
			  INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",
             INITP_00 => X"65AA996AA65AA994952D2DCB72DED2E0D5DE0DD5D080D0D5488DD63A80800008",
             INITP_01 => X"48D5DD5DD5DB7B7996AA65AA996AB0003000300020000200003577577576DEDE",
             INITP_02 => X"DD5DD5DB7B7996AA65AA996AB000D548D5DD5DD5DB7B7996AA65AA996AB000D5",
             INITP_03 => X"B7B7996AA65AA996ADB6DB6DD548D5DD5DD5DB7B7996AA65AA996AB000D548D5",
             INITP_04 => X"5DD5DB7B7996AA65AA996B5523577577576DEDE65AA996AA65AD548D5DD5DD5D",
             INITP_05 => X"00000000000000000000000000000000000000000000000000000000D548D5DD",
             INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
             INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000")
  --synthesis translate_on
port map(    DIA => "0000000000000000",
              DIPA => "00",
               ENA => '1',
               WEA => '0',
              SSRA => '0',
              CLKA => clk,
             ADDRA => addressA,
               DOA => instructionA(15 downto 0),
              DOPA => instructionA(17 downto 16),
      DIB => "0000000000000000",
              DIPB => "00",
               ENB => '1',
               WEB => '0',
              SSRB => '0',
              CLKB => clk,
             ADDRB => addressB,
               DOB => instructionB(15 downto 0),
              DOPB => instructionB(17 downto 16));  
--
end low_level_definition;
--
------------------------------------------------------------------------------------
--
-- END OF FILE lcd_prg.vhd
--
------------------------------------------------------------------------------------

